* C:\Users\shuof\PycharmProjects\capstone\test_data\MC1552G.asc
R1 VCC N002 9.0k
R2 VCC N003 5.0k
R3 VCC N001 500
Q4 VCC N001 Output 0 2N3904
Q3 N001 N003 N005 0 2N3904
Q2 N003 N002 0 0 2N3904
C1 N002 N003 3.0p
Q1 N002 Input N004 0 2N3904
R4 N005 N004 1.0k
R5 N004 0 150
C2 N005 N004 2.0p
R6 N005 0 80
R8 Output 0 3.0k
RK Output N006 6.0k
R7 0 Input 12k
Q6 0 N006 0 0 2N3904
Q8 Output N006 0 0 2N3904
D1_Q5 VCC Output D
D2_Q7 N006 0 D
R9 0 Gain_Select_Input_1 130
V1 VCC 0 6
C3 VCC 0 0.1u
R11 Vi 0 50
C4 Input Vi 0.01u
C5 0 0 5.0u
C6 Vo Output 0.1u
R12 Vo 0 1.0k
V2 Vi 0 AC 1
.model D D
.lib C:\Users\shuof\Documents\LTspiceXVII\lib\cmp\standard.dio
.model NPN NPN
.model PNP PNP
.lib C:\Users\shuof\Documents\LTspiceXVII\lib\cmp\standard.bjt
.op
.backanno
.end
