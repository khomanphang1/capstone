* C:\Users\shuof\PycharmProjects\capstone\test_data\2N3904_cascode.asc
V1 VCC 0 20
R1 VCC VB1 51k
R4 VCC VC1 5.5k
R2 VB1 VB2 3k
R3 VB2 0 5k
Q1 VC1 VB1 N001 0 2N3904
Q2 N001 VB2 N003 0 2N3904
R5 N003 N004 97.5
R6 N004 0 402.5
C4 N004 0 10u
C2 VB1 0 1u
C1 VB2 N002 1u
Rs N002 Vin 1k
V2 Vin 0 SINE(0 1 100K)
C3 VC1 Vout 1u
RL 0 Vout 100K
.model NPN NPN
.model PNP PNP
.lib C:\Users\shuof\Documents\LTspiceXVII\lib\cmp\standard.bjt
.op
.backanno
.end
