* C:\Users\shuof\PycharmProjects\capstone\test_data\ideal_common_source.asc
RS Vs 0 5k
RD 0 Vo 30k
Ro Vo Vs 200k
G1 Vo Vs Vs Vs 10e-3
Vi Vs 0 V
.backanno
.end
