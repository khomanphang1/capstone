Version 4
SHEET 1 1264 680
WIRE 240 -48 240 -112
WIRE 240 48 240 32
WIRE 352 48 240 48
WIRE 400 48 352 48
WIRE 464 48 400 48
WIRE 576 48 544 48
WIRE 304 96 240 96
WIRE 192 128 64 128
WIRE 304 144 304 96
WIRE 304 144 240 144
WIRE 400 160 400 48
WIRE 576 160 576 48
WIRE 240 176 240 144
WIRE 304 224 240 224
WIRE 80 256 64 256
WIRE 192 256 160 256
WIRE 240 272 240 256
WIRE 304 272 304 224
WIRE 304 272 240 272
WIRE 400 304 400 224
WIRE 576 304 576 240
WIRE 240 320 240 272
WIRE 400 320 400 304
FLAG 400 304 0
FLAG 240 320 0
FLAG 240 -112 0
FLAG 352 48 Vout
IOPIN 352 48 Out
FLAG -288 256 0
FLAG -304 16 0
FLAG -304 -64 Vbias
FLAG -288 176 Vin
FLAG 64 128 Vbias
FLAG 64 256 Vin
FLAG 576 304 0
SYMBOL current 240 -48 R0
SYMATTR InstName Ibias1
SYMATTR Value 0.25mA
SYMBOL cap 384 160 R0
SYMATTR InstName C_L
SYMATTR Value 4e-12
SYMBOL res 176 240 R90
WINDOW 0 0 56 VBottom 2
WINDOW 3 32 56 VTop 2
SYMATTR InstName Rs1
SYMATTR Value 10k
SYMBOL voltage -288 160 R0
SYMATTR InstName Vin1
SYMATTR Value 1
SYMATTR Value2 AC 1
SYMBOL voltage -304 -80 R0
SYMATTR InstName Vbias1
SYMATTR Value 2
SYMBOL nmos4 192 48 R0
SYMATTR InstName M1
SYMATTR Value NMOS0P5
SYMATTR Value2 l=10u w=1000u
SYMBOL nmos4 192 176 R0
SYMATTR InstName M2
SYMATTR Value NMOS0P5
SYMATTR Value2 l=10u w=1000u
SYMBOL res 560 32 R90
WINDOW 0 0 56 VBottom 2
WINDOW 3 32 56 VTop 2
SYMATTR InstName R_L
SYMATTR Value 1k
SYMBOL voltage 576 144 R0
SYMATTR InstName Vout_bias
SYMATTR Value 2V
TEXT 488 -200 Left 2 ;Hanspeter Schmid circuit
TEXT 504 -96 Left 2 !.model	NMOS0P5	NMOS(Level=1 VTO=0.5 KP= 20u LAMBDA=0.04)
TEXT 768 80 Left 2 ;HS values\ngm_1 = 1e-3\ngm_2 = 1e-3\nG_s = 1e-3\ng_ds1 = 1e-5\ng_ds2 = 1e-5\nC_L = 4e-12\nC_gs1 = 1e-13\nC_gs2 = 1e-13\nC-gd1 = 5e-15\nC_gd2 = 5e-15
TEXT 480 416 Left 2 !.op
