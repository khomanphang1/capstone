* C:\Users\shuof\PycharmProjects\capstone\test_data\ideal_common_source.asc
RS Vs 0 5k
RD 0 Vo 30k
Ro Vo Vs 200k
G1 Vo Vs Vg Vs 10e-3
Vi Vg 0 1
.backanno
.end
