* C:\Users\shuof\PycharmProjects\capstone\test_data\2N3904_common_emitter.asc
Q1 VC VB VE 0 2N3904
RC VCC VC 10k
RE VE 0 1k
R1 VCC VB 100k
R2 VB 0 100k
C1 VB Vin 16u
C2 N001 VE 3m
C3 VC Vout 160n
R3 N001 0 6
V1 VCC 0 9
V2 Vin 0 SINE(0 10m 1k)
RL Vout 0 100k
.model NPN NPN
.model PNP PNP
.lib C:\Users\shuof\Documents\LTspiceXVII\lib\cmp\standard.bjt
.op
.backanno
.end
