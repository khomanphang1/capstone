* C:\Users\shuof\PycharmProjects\capstone\test_data\transresistance.asc
Is 0 Vn 1m
Rid 0 Vn 100k
RF Vn Vo 10k
E1 Voc 0 0 Vn 100
Ro Vo Voc 1k
.backanno
.end
