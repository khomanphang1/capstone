* C:\Users\shuof\PycharmProjects\capstone\test_data\transresistance.asc
E1 Voc 0 0 Vp 100
Ro Voc Vo 200k
Rid Vp 0 10k
RF Vo Vp 5k
Is 0 Vp I
.backanno
.end
